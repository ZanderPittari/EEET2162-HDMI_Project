// D-Type Flip Flop

module dtype (
	input d;				// Data
	input clr_n;		// Clear
	input clk;			// Clock
	
	output q;			// Output
	output ld;			// Load

);

always @(clk)
	begin
		
	end

endmodule
